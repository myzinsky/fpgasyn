--
-- ROMs Using Block RAM Resources.
-- VHDL code for a ROM with registered output (template 1)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
entity blockrom is
    port ( clk   : in std_logic;
           en    : in std_logic;
           addr  : in std_logic_vector(7 downto 0);
           rec   : out integer range 0 to 909091;
           saw_n : out integer range 0 to 1818181;
           saw_m : out integer range 0 to 1417);
end blockrom;
architecture syn of blockrom is
    type rom_type is array (0 to 87) of integer range 0 to 1818181;
    signal ROM1 : rom_type:= (
				5919   , 6313   , 6576   , 7102   , 7398   , 7891   , 8523   , 8878  ,
				9470   , 9864   , 10522  , 11364  , 11837  , 12626  , 13152  , 14205 ,
				14796  , 15783  , 17045  , 17756  , 18939  , 19729  , 21044  , 22727 ,
				23674  , 25253  , 26305  , 28409  , 29593  , 31566  , 34091  , 35511 ,
				37879  , 39457  , 42088  , 45455  , 47348  , 50505  , 52609  , 56818 ,
				59186  , 63131  , 68182  , 71023  , 75758  , 78914  , 84175  , 90909 ,
				94697  , 101010 , 105219 , 113636 , 118371 , 126263 , 136364 , 142045,
				151515 , 157828 , 168350 , 181818 , 189394 , 202020 , 210438 , 227273,
				236742 , 252525 , 272727 , 284091 , 303030 , 315657 , 336700 , 363636,
				378788 , 404040 , 420875 , 454545 , 473485 , 505051 , 545455 , 568182,
				606061 , 631313 , 673401 , 727273 , 757576 , 808081 , 841751 , 909091
			    );

    signal ROM2 : rom_type:= (
				11837   , 12626   , 13152   , 14204   , 14796   , 15782    , 17045    , 17755   , 
				18939   , 19728   , 21043   , 22727   , 23674   , 25252    , 26304    , 28409   , 
				29592   , 31565   , 34090   , 35511   , 37878   , 39457    , 42087    , 45454   , 
				47348   , 50505   , 52609   , 56818   , 59185   , 63131    , 68181    , 71022   , 
				75757   , 78914   , 84175   , 90909   , 94696   , 101010   , 105218   , 113636  , 
				118371  , 126262  , 136363  , 142045  , 151515  , 157828   , 168350   , 181818  ,
				189393  , 202020  , 210437  , 227272  , 236742  , 252525   , 272727   , 284090  ,
				303030  , 315656  , 336700  , 363636  , 378787  , 404040   , 420875   , 454545  , 
				473484  , 505050  , 545454  , 568181  , 606060  , 631313   , 673400   , 727272  , 
				757575  , 808080  , 841750  , 909090  , 946969  , 1010101  , 1090909  , 1136363 , 
				1212121 , 1262626 , 1346801 , 1454545 , 1515151 , 1616161  , 1683501  , 1818181  
			    );

    signal ROM3 : rom_type:= (
				1417	, 1328	, 1275	, 1181	, 1133	, 1063	, 984	, 944	, 
				885	, 850	, 797	, 738	, 708	, 664	, 637	, 590	, 
				566	, 531	, 492	, 472	, 442	, 425	, 398	, 369	, 
				354	, 332	, 318	, 295	, 283	, 265	, 246	, 236	, 
				221	, 212	, 199	, 184	, 177	, 166	, 159	, 147	, 
				141	, 132	, 123	, 118	, 110	, 106	, 99	, 92	, 
				88	, 83	, 79	, 73	, 70	, 66	, 61	, 59	, 
				55	, 53	, 49	, 46	, 44	, 41	, 39	, 36	, 
				35	, 33	, 30	, 29	, 27	, 26	, 24	, 23	, 
				22	, 20	, 19	, 18	, 17	, 16	, 15	, 14	, 
				13	, 13	, 12	, 11	, 11	, 10	, 9	, 9
			    );

    signal real_addr : std_logic_vector(7 downto 0);

    signal data2 : integer range 0 to 909091;

begin

	real_addr <= X"6C" - addr ;

    process (clk)
    begin
        if (clk'event and clk = '1') then
             if (en = '1') then
                  rec   <= ROM1(conv_integer(real_addr));
                  saw_n <= ROM2(conv_integer(real_addr));
                  saw_m <= ROM3(conv_integer(real_addr));
             end if;
         end if;
    end process;
end syn;
